/* verilator lint_off MULTITOP */
module Hazard_detection_unit (
/* verilator lint_on MULTITOP */
	//inputs
//	input logic [1:0] WBSel_EX,
/* verilator lint_off UNUSED */
	input logic PCSel_EX,th1,
	input logic [4:0] rd_EX,rs1_ID,rs2_ID,rd_MEM,rs1_EX,rs2_EX,rd_WB,
	input logic [6:0] op_ex,op_id,
	input logic [31:0] pc_ID,alu,pc_EX,
/* verilator lint_on UNUSED */
	//outputs
	output logic stall_PC,stall_ID,flush_ID_EX,flush_IF_ID,
	output logic  comp_o,
	output logic  [31:0] PC_jump_EX
);
logic [31:0] temp;
always_comb begin
	case(PCSel_EX)
		1'b1: temp = alu;
		1'b0: temp = pc_EX + 32'h4;
		default: temp = 32'b0;
	endcase
//lw stall
	if(((rs1_ID == rd_EX) || (rs2_ID == rd_EX)) && (op_ex == 7'b0000011)) begin
		stall_PC = 1'b1;
		stall_ID = 1'b1;
		flush_IF_ID = 1'b0;
		flush_ID_EX  = 1'b1; 
	end else begin
		stall_PC = 1'b0;
		stall_ID = 1'b0;
		flush_IF_ID = 1'b0;
		flush_ID_EX  = 1'b0; 		
	end
// stall branch sat nhau
	if(th1)begin
		stall_PC = 1'b1;
		stall_ID = 1'b1;
		flush_IF_ID = 1'b0;
		flush_ID_EX = 1'b1;
	end else begin
		stall_PC = 1'b0;
		stall_ID = 1'b0;
		flush_IF_ID = 1'b0;
		flush_ID_EX = 1'b0;			
	end
//compare de fix		
	if(op_ex[6:4] != 3'b110)  begin
		comp_o = 1'b0;
	    flush_ID_EX = 1'b0;
		flush_IF_ID = 1'b0;	
	end else
		if(temp == pc_ID) begin
		comp_o = 1'b0;
	    flush_ID_EX = 1'b0;
		flush_IF_ID = 1'b0;
	end else begin
		comp_o = 1'b1;
		flush_ID_EX = 1'b1;
		flush_IF_ID = 1'b1;
	end

PC_jump_EX = temp; 
	
end
endmodule
